library verilog;
use verilog.vl_types.all;
entity testLab_vlg_vec_tst is
end testLab_vlg_vec_tst;
